library verilog;
use verilog.vl_types.all;
entity delay_vlg_check_tst is
    port(
        b               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end delay_vlg_check_tst;
