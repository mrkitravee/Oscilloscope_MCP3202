library verilog;
use verilog.vl_types.all;
entity Ossiloscope_MCP3202_vlg_vec_tst is
end Ossiloscope_MCP3202_vlg_vec_tst;
