library verilog;
use verilog.vl_types.all;
entity delay_vlg_vec_tst is
end delay_vlg_vec_tst;
