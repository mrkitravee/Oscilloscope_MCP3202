library verilog;
use verilog.vl_types.all;
entity Sending_WDATA_vlg_vec_tst is
end Sending_WDATA_vlg_vec_tst;
